module FFT_stage3(
input wire CLK,nRESET,stage2_done,
input wire signed [11:0] x_stage2_real [0:7],   //7 integer   5 fraction
input wire signed [11:0] x_stage2_image [0:7],   //7 integer   5 fraction
output reg signed [11:0] x_stage3_real [0:7],   //8 integer   4 fraction
output reg signed [11:0] x_stage3_image [0:7],   //8 integer   4 fraction
output reg stage3_done
);


reg signed [12:0] x_stage2_real_ex [0:7];
reg signed [12:0] x_stage2_image_ex [0:7];

always@(posedge CLK or negedge nRESET)
begin
    if(stage3_done)
       stage3_done <= 1'b0;

    if(!nRESET)
    begin
        stage3_done<=1'b0;
        for(int i=0; i<8; i=i+1)
        begin
            x_stage3_real[i] <=12'sd0;
            x_stage3_image[i] <=12'sd0;
        end
    end
    else if(stage2_done) begin

    for(int i=0; i<8 ; i=i+1)
    begin
            x_stage2_real_ex[i]= {x_stage2_real[i][11], x_stage2_real[i]};
            x_stage2_image_ex[i]= {x_stage2_image[i][11], x_stage2_image[i]};
    end

    x_stage3_real[0] <= ((x_stage2_real_ex[0] + x_stage2_real_ex[1]) >> 1);
    x_stage3_image[0] <= ((x_stage2_image_ex[0] + x_stage2_image_ex[1]) >> 1);

    x_stage3_real[2] <= ((x_stage2_real_ex[2] + x_stage2_real_ex[3]) >> 1);
    x_stage3_image[2] <= ((x_stage2_image_ex[2] + x_stage2_image_ex[3]) >> 1);

    x_stage3_real[4] <= ((x_stage2_real_ex[4] + x_stage2_real_ex[5]) >> 1);
    x_stage3_image[4] <= ((x_stage2_image_ex[4] + x_stage2_image_ex[5]) >> 1);

    x_stage3_real[6] <= ((x_stage2_real_ex[6] + x_stage2_real_ex[7]) >> 1);
    x_stage3_image[6] <= ((x_stage2_image_ex[6] + x_stage2_image_ex[7]) >> 1);




    x_stage3_real[1] <= ((x_stage2_real_ex[0] - x_stage2_real_ex[1]) >> 1);
    x_stage3_image[1] <= ((x_stage2_image_ex[0] - x_stage2_image_ex[1]) >> 1); 

    x_stage3_real[3] <= ((x_stage2_real_ex[2] - x_stage2_real_ex[3]) >> 1);
    x_stage3_image[3] <= ((x_stage2_image_ex[2] - x_stage2_image_ex[3]) >> 1);

    x_stage3_real[5] <= ((x_stage2_real_ex[4] - x_stage2_real_ex[5]) >> 1);
    x_stage3_image[5] <= ((x_stage2_image_ex[4] - x_stage2_image_ex[5]) >> 1);

    x_stage3_real[7] <= ((x_stage2_real_ex[6] - x_stage2_real_ex[7]) >> 1);
    x_stage3_image[7] <= ((x_stage2_image_ex[6] - x_stage2_image_ex[7]) >> 1);


    stage3_done<=1'b1;              
    end
end
endmodule